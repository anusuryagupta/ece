----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/18/2025 09:03:12 AM
-- Design Name: 
-- Module Name: lab9 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library xil_defaultlib;
use xil_defaultlib.all;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity fourbitregister is
    Port (clk : in STD_LOGIC;
          d : in STD_LOGIC_VECTOR(3 downto 0);
          q : out STD_LOGIC_VECTOR(3 downto 0));
end fourbitregister;

architecture Behavioral of fourbitregister is

begin
    process(clk)
        begin
        if rising_edge(clk) then
            q <= d;
        end if;
    end process;
end Behavioral;
